###############################################################################
#TSMC Library/IP Product
#Filename: tpzn65lpgv2od3_9lm.lef
#Technology: CLN65LP
#Product Type: Standard I/O
#Product Name: tpzn65lpgv2od3
#Version: 200b
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.005 BY 190.000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 190.000 BY 190.000 ;
END corner

MACRO PCI33DGZ
    CLASS PAD ;
    FOREIGN PCI33DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PCI33DGZ

MACRO PCI33SDGZ
    CLASS PAD ;
    FOREIGN PCI33SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PCI33SDGZ

MACRO PCI66DGZ
    CLASS PAD ;
    FOREIGN PCI66DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PCI66DGZ

MACRO PCI66SDGZ
    CLASS PAD ;
    FOREIGN PCI66SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PCI66SDGZ

MACRO PCLAMP1ANA
    CLASS BLOCK ;
    FOREIGN PCLAMP1ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 106.605 BY 65.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        DIRECTION INOUT ;
        PORT
        LAYER M3 ;
        RECT  55.910 0.000 57.410 9.000 ;
        RECT  55.910 56.000 57.410 65.000 ;
        RECT  52.480 0.000 54.320 9.000 ;
        RECT  52.480 56.000 54.320 65.000 ;
        RECT  46.350 0.000 50.030 9.000 ;
        RECT  46.350 56.000 50.030 65.000 ;
        RECT  39.680 0.000 43.360 9.000 ;
        RECT  39.680 56.000 43.360 65.000 ;
        RECT  33.550 0.000 37.230 9.000 ;
        RECT  33.550 56.000 37.230 65.000 ;
        RECT  27.890 0.000 31.100 9.000 ;
        RECT  27.890 56.000 31.100 65.000 ;
        RECT  21.760 0.000 25.440 9.000 ;
        RECT  21.760 56.000 25.440 65.000 ;
        RECT  15.090 0.000 19.810 9.000 ;
        RECT  15.090 56.000 19.810 65.000 ;
        RECT  8.960 0.000 12.640 9.000 ;
        RECT  8.960 56.000 12.640 65.000 ;
        RECT  1.500 0.000 6.510 2.000 ;
        RECT  1.500 13.875 6.510 18.375 ;
        RECT  1.500 30.250 6.510 34.750 ;
        RECT  1.500 46.625 6.510 51.125 ;
        RECT  1.500 63.000 6.510 65.000 ;
        END
    END VSSESD
    PIN VDDESD
        DIRECTION INOUT ;
        PORT
        LAYER M3 ;
        RECT  96.105 0.000 105.105 2.000 ;
        RECT  96.105 13.875 105.105 18.375 ;
        RECT  96.105 30.250 105.105 34.750 ;
        RECT  96.105 46.625 105.105 51.125 ;
        RECT  96.105 63.000 105.105 65.000 ;
        RECT  91.105 0.000 96.105 9.000 ;
        RECT  91.105 56.000 96.105 65.000 ;
        RECT  82.105 0.000 87.105 9.000 ;
        RECT  82.105 56.000 87.105 65.000 ;
        RECT  73.105 0.000 78.105 9.000 ;
        RECT  73.105 56.000 78.105 65.000 ;
        RECT  64.105 0.000 69.105 9.000 ;
        RECT  64.105 56.000 69.105 65.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 106.605 65.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 106.605 65.000 ;
        LAYER VIA2 ;
        RECT  96.105 0.000 105.105 2.000 ;
        RECT  96.105 63.000 105.105 65.000 ;
        RECT  91.105 0.000 96.105 9.000 ;
        RECT  91.105 56.000 96.105 65.000 ;
        RECT  82.105 0.000 87.105 9.000 ;
        RECT  82.105 56.000 87.105 65.000 ;
        RECT  73.105 0.000 78.105 9.000 ;
        RECT  73.105 56.000 78.105 65.000 ;
        RECT  64.105 0.000 69.105 9.000 ;
        RECT  64.105 56.000 69.105 65.000 ;
        RECT  55.910 0.000 57.410 9.000 ;
        RECT  55.910 56.000 57.410 65.000 ;
        RECT  52.480 0.000 54.320 9.000 ;
        RECT  52.480 56.000 54.320 65.000 ;
        RECT  46.350 0.000 50.030 9.000 ;
        RECT  46.350 56.000 50.030 65.000 ;
        RECT  39.680 0.000 43.360 9.000 ;
        RECT  39.680 56.000 43.360 65.000 ;
        RECT  33.550 0.000 37.230 9.000 ;
        RECT  33.550 56.000 37.230 65.000 ;
        RECT  27.890 0.000 31.100 9.000 ;
        RECT  27.890 56.000 31.100 65.000 ;
        RECT  21.760 0.000 25.440 9.000 ;
        RECT  21.760 56.000 25.440 65.000 ;
        RECT  15.090 0.000 19.810 9.000 ;
        RECT  15.090 56.000 19.810 65.000 ;
        RECT  8.960 0.000 12.640 9.000 ;
        RECT  8.960 56.000 12.640 65.000 ;
        LAYER M3 ;
        RECT  105.605 0.000 106.605 65.000 ;
        RECT  97.605 2.500 105.605 62.500 ;
        RECT  89.605 10.500 97.605 54.500 ;
        RECT  88.605 0.000 89.605 65.000 ;
        RECT  80.605 10.500 88.605 54.500 ;
        RECT  79.605 0.000 80.605 65.000 ;
        RECT  71.605 10.500 79.605 54.500 ;
        RECT  70.605 0.000 71.605 65.000 ;
        RECT  62.605 10.500 70.605 54.500 ;
        RECT  57.570 0.000 62.605 65.000 ;
        RECT  55.750 9.160 57.570 55.840 ;
        RECT  54.820 0.000 55.750 65.000 ;
        RECT  51.980 9.500 54.820 55.500 ;
        RECT  50.530 0.000 51.980 65.000 ;
        RECT  45.850 9.500 50.530 55.500 ;
        RECT  43.860 0.000 45.850 65.000 ;
        RECT  39.180 9.500 43.860 55.500 ;
        RECT  37.730 0.000 39.180 65.000 ;
        RECT  33.050 9.500 37.730 55.500 ;
        RECT  31.600 0.000 33.050 65.000 ;
        RECT  27.390 9.500 31.600 55.500 ;
        RECT  25.940 0.000 27.390 65.000 ;
        RECT  21.310 9.500 25.940 55.500 ;
        RECT  13.590 10.500 21.310 54.500 ;
        RECT  13.140 0.000 13.590 65.000 ;
        RECT  8.460 9.500 13.140 55.500 ;
        RECT  7.010 0.000 8.460 65.000 ;
        RECT  1.000 2.500 7.010 62.500 ;
        RECT  0.000 0.000 1.000 65.000 ;
    END
END PCLAMP1ANA

MACRO PCLAMP2ANA
    CLASS BLOCK ;
    FOREIGN PCLAMP2ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 106.605 BY 65.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        DIRECTION INOUT ;
        PORT
        LAYER M3 ;
        RECT  55.910 0.000 57.410 9.000 ;
        RECT  55.910 56.000 57.410 65.000 ;
        RECT  52.480 0.000 54.320 9.000 ;
        RECT  52.480 56.000 54.320 65.000 ;
        RECT  46.350 0.000 50.030 9.000 ;
        RECT  46.350 56.000 50.030 65.000 ;
        RECT  39.680 0.000 43.360 9.000 ;
        RECT  39.680 56.000 43.360 65.000 ;
        RECT  33.550 0.000 37.230 9.000 ;
        RECT  33.550 56.000 37.230 65.000 ;
        RECT  27.890 0.000 31.100 9.000 ;
        RECT  27.890 56.000 31.100 65.000 ;
        RECT  21.760 0.000 25.440 9.000 ;
        RECT  21.760 56.000 25.440 65.000 ;
        RECT  15.090 0.000 19.810 9.000 ;
        RECT  15.090 56.000 19.810 65.000 ;
        RECT  8.960 0.000 12.640 9.000 ;
        RECT  8.960 56.000 12.640 65.000 ;
        RECT  1.500 0.000 6.510 2.000 ;
        RECT  1.500 13.875 6.510 18.375 ;
        RECT  1.500 30.250 6.510 34.750 ;
        RECT  1.500 46.625 6.510 51.125 ;
        RECT  1.500 63.000 6.510 65.000 ;
        END
    END VSSESD
    PIN VDDESD
        DIRECTION INOUT ;
        PORT
        LAYER M3 ;
        RECT  96.105 0.000 105.105 2.000 ;
        RECT  96.105 13.875 105.105 18.375 ;
        RECT  96.105 30.250 105.105 34.750 ;
        RECT  96.105 46.625 105.105 51.125 ;
        RECT  96.105 63.000 105.105 65.000 ;
        RECT  91.105 0.000 96.105 9.000 ;
        RECT  91.105 56.000 96.105 65.000 ;
        RECT  82.105 0.000 87.105 9.000 ;
        RECT  82.105 56.000 87.105 65.000 ;
        RECT  73.105 0.000 78.105 9.000 ;
        RECT  73.105 56.000 78.105 65.000 ;
        RECT  64.105 0.000 69.105 9.000 ;
        RECT  64.105 56.000 69.105 65.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 106.605 65.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 106.605 65.000 ;
        LAYER VIA2 ;
        RECT  96.105 0.000 105.105 2.000 ;
        RECT  96.105 63.000 105.105 65.000 ;
        RECT  91.105 0.000 96.105 9.000 ;
        RECT  91.105 56.000 96.105 65.000 ;
        RECT  82.105 0.000 87.105 9.000 ;
        RECT  82.105 56.000 87.105 65.000 ;
        RECT  73.105 0.000 78.105 9.000 ;
        RECT  73.105 56.000 78.105 65.000 ;
        RECT  64.105 0.000 69.105 9.000 ;
        RECT  64.105 56.000 69.105 65.000 ;
        RECT  55.910 0.000 57.410 9.000 ;
        RECT  55.910 56.000 57.410 65.000 ;
        RECT  52.480 0.000 54.320 9.000 ;
        RECT  52.480 56.000 54.320 65.000 ;
        RECT  46.350 0.000 50.030 9.000 ;
        RECT  46.350 56.000 50.030 65.000 ;
        RECT  39.680 0.000 43.360 9.000 ;
        RECT  39.680 56.000 43.360 65.000 ;
        RECT  33.550 0.000 37.230 9.000 ;
        RECT  33.550 56.000 37.230 65.000 ;
        RECT  27.890 0.000 31.100 9.000 ;
        RECT  27.890 56.000 31.100 65.000 ;
        RECT  21.760 0.000 25.440 9.000 ;
        RECT  21.760 56.000 25.440 65.000 ;
        RECT  15.090 0.000 19.810 9.000 ;
        RECT  15.090 56.000 19.810 65.000 ;
        RECT  8.960 0.000 12.640 9.000 ;
        RECT  8.960 56.000 12.640 65.000 ;
        LAYER M3 ;
        RECT  105.605 0.000 106.605 65.000 ;
        RECT  97.605 2.500 105.605 62.500 ;
        RECT  89.605 10.500 97.605 54.500 ;
        RECT  88.605 0.000 89.605 65.000 ;
        RECT  80.605 10.500 88.605 54.500 ;
        RECT  79.605 0.000 80.605 65.000 ;
        RECT  71.605 10.500 79.605 54.500 ;
        RECT  70.605 0.000 71.605 65.000 ;
        RECT  62.605 10.500 70.605 54.500 ;
        RECT  57.570 0.000 62.605 65.000 ;
        RECT  55.750 9.160 57.570 55.840 ;
        RECT  54.820 0.000 55.750 65.000 ;
        RECT  51.980 9.500 54.820 55.500 ;
        RECT  50.530 0.000 51.980 65.000 ;
        RECT  45.850 9.500 50.530 55.500 ;
        RECT  43.860 0.000 45.850 65.000 ;
        RECT  39.180 9.500 43.860 55.500 ;
        RECT  37.730 0.000 39.180 65.000 ;
        RECT  33.050 9.500 37.730 55.500 ;
        RECT  31.600 0.000 33.050 65.000 ;
        RECT  27.390 9.500 31.600 55.500 ;
        RECT  25.940 0.000 27.390 65.000 ;
        RECT  21.310 9.500 25.940 55.500 ;
        RECT  13.590 10.500 21.310 54.500 ;
        RECT  13.140 0.000 13.590 65.000 ;
        RECT  8.460 9.500 13.140 55.500 ;
        RECT  7.010 0.000 8.460 65.000 ;
        RECT  1.000 2.500 7.010 62.500 ;
        RECT  0.000 0.000 1.000 65.000 ;
    END
END PCLAMP2ANA

MACRO PCORNER
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNER 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 190.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE corner ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 190.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 190.000 190.000 ;
    END
END PCORNER

MACRO PDB02DGZ
    CLASS PAD ;
    FOREIGN PDB02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB02DGZ

MACRO PDB02SDGZ
    CLASS PAD ;
    FOREIGN PDB02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB02SDGZ

MACRO PDB04DGZ
    CLASS PAD ;
    FOREIGN PDB04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB04DGZ

MACRO PDB04SDGZ
    CLASS PAD ;
    FOREIGN PDB04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB04SDGZ

MACRO PDB08DGZ
    CLASS PAD ;
    FOREIGN PDB08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB08DGZ

MACRO PDB08SDGZ
    CLASS PAD ;
    FOREIGN PDB08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB08SDGZ

MACRO PDB12DGZ
    CLASS PAD ;
    FOREIGN PDB12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB12DGZ

MACRO PDB12SDGZ
    CLASS PAD ;
    FOREIGN PDB12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB12SDGZ

MACRO PDB16DGZ
    CLASS PAD ;
    FOREIGN PDB16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB16DGZ

MACRO PDB16SDGZ
    CLASS PAD ;
    FOREIGN PDB16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB16SDGZ

MACRO PDB24DGZ
    CLASS PAD ;
    FOREIGN PDB24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB24DGZ

MACRO PDB24SDGZ
    CLASS PAD ;
    FOREIGN PDB24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDB24SDGZ

MACRO PDD02DGZ
    CLASS PAD ;
    FOREIGN PDD02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD02DGZ

MACRO PDD02SDGZ
    CLASS PAD ;
    FOREIGN PDD02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD02SDGZ

MACRO PDD04DGZ
    CLASS PAD ;
    FOREIGN PDD04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD04DGZ

MACRO PDD04SDGZ
    CLASS PAD ;
    FOREIGN PDD04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD04SDGZ

MACRO PDD08DGZ
    CLASS PAD ;
    FOREIGN PDD08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD08DGZ

MACRO PDD08SDGZ
    CLASS PAD ;
    FOREIGN PDD08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD08SDGZ

MACRO PDD12DGZ
    CLASS PAD ;
    FOREIGN PDD12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD12DGZ

MACRO PDD12SDGZ
    CLASS PAD ;
    FOREIGN PDD12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD12SDGZ

MACRO PDD16DGZ
    CLASS PAD ;
    FOREIGN PDD16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD16DGZ

MACRO PDD16SDGZ
    CLASS PAD ;
    FOREIGN PDD16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD16SDGZ

MACRO PDD24DGZ
    CLASS PAD ;
    FOREIGN PDD24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD24DGZ

MACRO PDD24SDGZ
    CLASS PAD ;
    FOREIGN PDD24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDD24SDGZ

MACRO PDDDGZ
    CLASS PAD ;
    FOREIGN PDDDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDDDGZ

MACRO PDDSDGZ
    CLASS PAD ;
    FOREIGN PDDSDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDDSDGZ

MACRO PDDW02DGZ
    CLASS PAD ;
    FOREIGN PDDW02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW02DGZ

MACRO PDDW04DGZ
    CLASS PAD ;
    FOREIGN PDDW04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW04DGZ

MACRO PDDW08DGZ
    CLASS PAD ;
    FOREIGN PDDW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW08DGZ

MACRO PDDW12DGZ
    CLASS PAD ;
    FOREIGN PDDW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW12DGZ

MACRO PDDW16DGZ
    CLASS PAD ;
    FOREIGN PDDW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW16DGZ

MACRO PDDW24DGZ
    CLASS PAD ;
    FOREIGN PDDW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDDW24DGZ

MACRO PDDWDGZ
    CLASS PAD ;
    FOREIGN PDDWDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  3.500 88.185 18.505 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDDWDGZ

MACRO PDIDGZ
    CLASS PAD ;
    FOREIGN PDIDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDIDGZ

MACRO PDISDGZ
    CLASS PAD ;
    FOREIGN PDISDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDISDGZ

MACRO PDO02CDG
    CLASS PAD ;
    FOREIGN PDO02CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO02CDG

MACRO PDO04CDG
    CLASS PAD ;
    FOREIGN PDO04CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO04CDG

MACRO PDO08CDG
    CLASS PAD ;
    FOREIGN PDO08CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO08CDG

MACRO PDO12CDG
    CLASS PAD ;
    FOREIGN PDO12CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO12CDG

MACRO PDO16CDG
    CLASS PAD ;
    FOREIGN PDO16CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO16CDG

MACRO PDO24CDG
    CLASS PAD ;
    FOREIGN PDO24CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDO24CDG

MACRO PDT02DGZ
    CLASS PAD ;
    FOREIGN PDT02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT02DGZ

MACRO PDT04DGZ
    CLASS PAD ;
    FOREIGN PDT04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT04DGZ

MACRO PDT08DGZ
    CLASS PAD ;
    FOREIGN PDT08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT08DGZ

MACRO PDT12DGZ
    CLASS PAD ;
    FOREIGN PDT12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT12DGZ

MACRO PDT16DGZ
    CLASS PAD ;
    FOREIGN PDT16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT16DGZ

MACRO PDT24DGZ
    CLASS PAD ;
    FOREIGN PDT24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDT24DGZ

MACRO PDU02DGZ
    CLASS PAD ;
    FOREIGN PDU02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU02DGZ

MACRO PDU02SDGZ
    CLASS PAD ;
    FOREIGN PDU02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU02SDGZ

MACRO PDU04DGZ
    CLASS PAD ;
    FOREIGN PDU04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU04DGZ

MACRO PDU04SDGZ
    CLASS PAD ;
    FOREIGN PDU04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU04SDGZ

MACRO PDU08DGZ
    CLASS PAD ;
    FOREIGN PDU08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU08DGZ

MACRO PDU08SDGZ
    CLASS PAD ;
    FOREIGN PDU08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU08SDGZ

MACRO PDU12DGZ
    CLASS PAD ;
    FOREIGN PDU12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU12DGZ

MACRO PDU12SDGZ
    CLASS PAD ;
    FOREIGN PDU12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU12SDGZ

MACRO PDU16DGZ
    CLASS PAD ;
    FOREIGN PDU16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU16DGZ

MACRO PDU16SDGZ
    CLASS PAD ;
    FOREIGN PDU16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU16SDGZ

MACRO PDU24DGZ
    CLASS PAD ;
    FOREIGN PDU24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU24DGZ

MACRO PDU24SDGZ
    CLASS PAD ;
    FOREIGN PDU24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDU24SDGZ

MACRO PDUDGZ
    CLASS PAD ;
    FOREIGN PDUDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDUDGZ

MACRO PDUSDGZ
    CLASS PAD ;
    FOREIGN PDUSDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  0.000 0.000 25.705 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  3.500 88.185 25.705 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDUSDGZ

MACRO PDUW02DGZ
    CLASS PAD ;
    FOREIGN PDUW02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW02DGZ

MACRO PDUW04DGZ
    CLASS PAD ;
    FOREIGN PDUW04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW04DGZ

MACRO PDUW08DGZ
    CLASS PAD ;
    FOREIGN PDUW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW08DGZ

MACRO PDUW12DGZ
    CLASS PAD ;
    FOREIGN PDUW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW12DGZ

MACRO PDUW16DGZ
    CLASS PAD ;
    FOREIGN PDUW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW16DGZ

MACRO PDUW24DGZ
    CLASS PAD ;
    FOREIGN PDUW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PDUW24DGZ

MACRO PDUWDGZ
    CLASS PAD ;
    FOREIGN PDUWDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  0.000 0.000 18.505 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  3.500 88.185 18.505 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDUWDGZ

MACRO PDXO01DG
    CLASS PAD ;
    FOREIGN PDXO01DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  38.500 88.185 49.910 190.000 ;
        RECT  26.500 0.000 38.500 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXO01DG

MACRO PDXO02DG
    CLASS PAD ;
    FOREIGN PDXO02DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  38.500 88.185 49.910 190.000 ;
        RECT  26.500 0.000 38.500 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXO02DG

MACRO PDXO03DG
    CLASS PAD ;
    FOREIGN PDXO03DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  0.000 0.000 49.910 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  38.500 88.185 49.910 190.000 ;
        RECT  26.500 0.000 38.500 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXO03DG

MACRO PDXOE1DG
    CLASS PAD ;
    FOREIGN PDXOE1DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M1 ;
        RECT  37.130 189.000 39.900 190.000 ;
        END
    END E
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  40.060 88.185 49.910 190.000 ;
        RECT  38.500 88.185 40.060 188.840 ;
        RECT  36.970 0.000 38.500 188.840 ;
        RECT  26.500 0.000 36.970 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXOE1DG

MACRO PDXOE2DG
    CLASS PAD ;
    FOREIGN PDXOE2DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M1 ;
        RECT  37.130 189.000 39.900 190.000 ;
        END
    END E
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  40.060 88.185 49.910 190.000 ;
        RECT  38.500 88.185 40.060 188.840 ;
        RECT  36.970 0.000 38.500 188.840 ;
        RECT  26.500 0.000 36.970 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXOE2DG

MACRO PDXOE3DG
    CLASS PAD ;
    FOREIGN PDXOE3DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M6 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M5 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M4 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M3 ;
        RECT  40.000 78.685 60.000 86.685 ;
        LAYER M2 ;
        RECT  47.210 0.750 52.790 1.750 ;
        RECT  40.000 78.685 60.000 86.685 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        LAYER M1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M1 ;
        RECT  37.130 189.000 39.900 190.000 ;
        END
    END E
    OBS
        LAYER M1 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA1 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M2 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA2 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M3 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA3 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M4 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA4 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M5 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA5 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M6 ;
        RECT  53.000 0.000 65.000 190.000 ;
        RECT  49.910 0.000 53.000 188.840 ;
        RECT  40.060 0.000 49.910 190.000 ;
        RECT  36.970 0.000 40.060 188.840 ;
        RECT  0.000 0.000 36.970 190.000 ;
        LAYER VIA6 ;
        RECT  50.070 189.000 52.840 190.000 ;
        RECT  37.130 189.000 39.900 190.000 ;
        LAYER M7 ;
        RECT  61.500 0.000 65.000 190.000 ;
        RECT  38.500 0.000 61.500 77.185 ;
        RECT  53.000 88.185 61.500 190.000 ;
        RECT  49.910 88.185 53.000 188.840 ;
        RECT  40.060 88.185 49.910 190.000 ;
        RECT  38.500 88.185 40.060 188.840 ;
        RECT  36.970 0.000 38.500 188.840 ;
        RECT  26.500 0.000 36.970 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PDXOE3DG

MACRO PFILLER0005
    CLASS PAD SPACER ;
    FOREIGN PFILLER0005 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.005 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.005 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.005 190.000 ;
    END
END PFILLER0005

MACRO PFILLER05
    CLASS PAD SPACER ;
    FOREIGN PFILLER05 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.500 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.500 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.500 190.000 ;
    END
END PFILLER05

MACRO PFILLER1
    CLASS PAD SPACER ;
    FOREIGN PFILLER1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 1.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 1.000 190.000 ;
    END
END PFILLER1

MACRO PFILLER10
    CLASS PAD SPACER ;
    FOREIGN PFILLER10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 10.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 10.000 190.000 ;
    END
END PFILLER10

MACRO PFILLER20
    CLASS PAD SPACER ;
    FOREIGN PFILLER20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 20.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 20.000 190.000 ;
    END
END PFILLER20

MACRO PFILLER5
    CLASS PAD SPACER ;
    FOREIGN PFILLER5 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 5.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 5.000 190.000 ;
    END
END PFILLER5

MACRO PRB08DGZ
    CLASS PAD ;
    FOREIGN PRB08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB08DGZ

MACRO PRB08SDGZ
    CLASS PAD ;
    FOREIGN PRB08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB08SDGZ

MACRO PRB12DGZ
    CLASS PAD ;
    FOREIGN PRB12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB12DGZ

MACRO PRB12SDGZ
    CLASS PAD ;
    FOREIGN PRB12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB12SDGZ

MACRO PRB16DGZ
    CLASS PAD ;
    FOREIGN PRB16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB16DGZ

MACRO PRB16SDGZ
    CLASS PAD ;
    FOREIGN PRB16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB16SDGZ

MACRO PRB24DGZ
    CLASS PAD ;
    FOREIGN PRB24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB24DGZ

MACRO PRB24SDGZ
    CLASS PAD ;
    FOREIGN PRB24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRB24SDGZ

MACRO PRCUT
    CLASS PAD ;
    FOREIGN PRCUT 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 30.000 190.000 ;
    END
END PRCUT

MACRO PRD08DGZ
    CLASS PAD ;
    FOREIGN PRD08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD08DGZ

MACRO PRD08SDGZ
    CLASS PAD ;
    FOREIGN PRD08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD08SDGZ

MACRO PRD12DGZ
    CLASS PAD ;
    FOREIGN PRD12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD12DGZ

MACRO PRD12SDGZ
    CLASS PAD ;
    FOREIGN PRD12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD12SDGZ

MACRO PRD16DGZ
    CLASS PAD ;
    FOREIGN PRD16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD16DGZ

MACRO PRD16SDGZ
    CLASS PAD ;
    FOREIGN PRD16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD16SDGZ

MACRO PRD24DGZ
    CLASS PAD ;
    FOREIGN PRD24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD24DGZ

MACRO PRD24SDGZ
    CLASS PAD ;
    FOREIGN PRD24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRD24SDGZ

MACRO PRDW08DGZ
    CLASS PAD ;
    FOREIGN PRDW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRDW08DGZ

MACRO PRDW12DGZ
    CLASS PAD ;
    FOREIGN PRDW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRDW12DGZ

MACRO PRDW16DGZ
    CLASS PAD ;
    FOREIGN PRDW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRDW16DGZ

MACRO PRDW24DGZ
    CLASS PAD ;
    FOREIGN PRDW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRDW24DGZ

MACRO PRO08CDG
    CLASS PAD ;
    FOREIGN PRO08CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRO08CDG

MACRO PRO12CDG
    CLASS PAD ;
    FOREIGN PRO12CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRO12CDG

MACRO PRO16CDG
    CLASS PAD ;
    FOREIGN PRO16CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRO16CDG

MACRO PRO24CDG
    CLASS PAD ;
    FOREIGN PRO24CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  3.930 0.000 30.000 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.930 88.185 26.500 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRO24CDG

MACRO PRT08DGZ
    CLASS PAD ;
    FOREIGN PRT08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRT08DGZ

MACRO PRT12DGZ
    CLASS PAD ;
    FOREIGN PRT12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRT12DGZ

MACRO PRT16DGZ
    CLASS PAD ;
    FOREIGN PRT16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRT16DGZ

MACRO PRT24DGZ
    CLASS PAD ;
    FOREIGN PRT24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    OBS
        LAYER M1 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  17.635 0.000 30.000 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  17.635 88.185 26.500 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRT24DGZ

MACRO PRU08DGZ
    CLASS PAD ;
    FOREIGN PRU08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU08DGZ

MACRO PRU08SDGZ
    CLASS PAD ;
    FOREIGN PRU08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU08SDGZ

MACRO PRU12DGZ
    CLASS PAD ;
    FOREIGN PRU12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU12DGZ

MACRO PRU12SDGZ
    CLASS PAD ;
    FOREIGN PRU12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU12SDGZ

MACRO PRU16DGZ
    CLASS PAD ;
    FOREIGN PRU16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU16DGZ

MACRO PRU16SDGZ
    CLASS PAD ;
    FOREIGN PRU16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU16SDGZ

MACRO PRU24DGZ
    CLASS PAD ;
    FOREIGN PRU24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU24DGZ

MACRO PRU24SDGZ
    CLASS PAD ;
    FOREIGN PRU24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  17.635 0.000 25.705 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  17.635 88.185 25.705 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRU24SDGZ

MACRO PRUW08DGZ
    CLASS PAD ;
    FOREIGN PRUW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRUW08DGZ

MACRO PRUW12DGZ
    CLASS PAD ;
    FOREIGN PRUW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRUW12DGZ

MACRO PRUW16DGZ
    CLASS PAD ;
    FOREIGN PRUW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRUW16DGZ

MACRO PRUW24DGZ
    CLASS PAD ;
    FOREIGN PRUW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M6 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M5 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M4 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M3 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M2 ;
        RECT  18.665 189.000 21.435 190.000 ;
        LAYER M1 ;
        RECT  18.665 189.000 21.435 190.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  12.210 0.750 17.790 1.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M6 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M5 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M4 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M3 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M2 ;
        RECT  14.705 189.000 17.475 190.000 ;
        LAYER M1 ;
        RECT  14.705 189.000 17.475 190.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M1 ;
        RECT  1.000 189.000 3.770 190.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        LAYER M1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        END
    END C
    OBS
        LAYER M1 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA1 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M2 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA2 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M3 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA3 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M4 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA4 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M5 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA5 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M6 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  25.705 0.000 28.795 188.840 ;
        RECT  21.595 0.000 25.705 190.000 ;
        RECT  18.505 0.000 21.595 188.840 ;
        RECT  17.635 0.000 18.505 190.000 ;
        RECT  14.545 0.000 17.635 188.840 ;
        RECT  3.930 0.000 14.545 190.000 ;
        RECT  0.840 0.000 3.930 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
        LAYER VIA6 ;
        RECT  25.865 189.000 28.635 190.000 ;
        RECT  18.665 189.000 21.435 190.000 ;
        RECT  14.705 189.000 17.475 190.000 ;
        RECT  1.000 189.000 3.770 190.000 ;
        LAYER M7 ;
        RECT  28.795 0.000 30.000 190.000 ;
        RECT  26.500 0.000 28.795 188.840 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  25.705 88.185 26.500 188.840 ;
        RECT  21.595 88.185 25.705 190.000 ;
        RECT  18.505 88.185 21.595 188.840 ;
        RECT  17.635 88.185 18.505 190.000 ;
        RECT  14.545 88.185 17.635 188.840 ;
        RECT  3.930 88.185 14.545 190.000 ;
        RECT  3.500 88.185 3.930 188.840 ;
        RECT  0.840 0.000 3.500 188.840 ;
        RECT  0.000 0.000 0.840 190.000 ;
    END
END PRUW24DGZ

MACRO PVDD1ANA
    CLASS PAD ;
    FOREIGN PVDD1ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AVDD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  15.630 0.750 16.690 1.365 ;
        RECT  5.000 78.685 25.000 86.680 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        LAYER M1 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  15.630 0.750 16.690 1.365 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  27.955 0.000 30.000 190.000 ;
        RECT  20.905 0.000 27.955 185.560 ;
        RECT  18.500 0.000 20.905 190.000 ;
        RECT  11.500 0.000 18.500 185.560 ;
        RECT  9.095 0.000 11.500 190.000 ;
        RECT  2.045 0.000 9.095 185.560 ;
        RECT  0.000 0.000 2.045 190.000 ;
        LAYER VIA1 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        LAYER M2 ;
        RECT  27.955 0.000 30.000 190.000 ;
        RECT  20.905 0.000 27.955 185.560 ;
        RECT  18.500 0.000 20.905 190.000 ;
        RECT  11.500 0.000 18.500 185.560 ;
        RECT  9.095 0.000 11.500 190.000 ;
        RECT  2.045 0.000 9.095 185.560 ;
        RECT  0.000 0.000 2.045 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVDD1ANA

MACRO PVDD1DGZ
    CLASS PAD ;
    FOREIGN PVDD1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  15.630 0.750 16.690 1.365 ;
        RECT  5.000 78.685 25.000 86.680 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        LAYER M1 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  15.630 0.750 16.690 1.365 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  27.955 0.000 30.000 190.000 ;
        RECT  20.905 0.000 27.955 185.560 ;
        RECT  18.500 0.000 20.905 190.000 ;
        RECT  11.500 0.000 18.500 185.560 ;
        RECT  9.095 0.000 11.500 190.000 ;
        RECT  2.045 0.000 9.095 185.560 ;
        RECT  0.000 0.000 2.045 190.000 ;
        LAYER VIA1 ;
        RECT  21.405 186.060 27.455 190.000 ;
        RECT  12.000 186.060 18.000 190.000 ;
        RECT  2.545 186.060 8.595 190.000 ;
        LAYER M2 ;
        RECT  27.955 0.000 30.000 190.000 ;
        RECT  20.905 0.000 27.955 185.560 ;
        RECT  18.500 0.000 20.905 190.000 ;
        RECT  11.500 0.000 18.500 185.560 ;
        RECT  9.095 0.000 11.500 190.000 ;
        RECT  2.045 0.000 9.095 185.560 ;
        RECT  0.000 0.000 2.045 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVDD1DGZ

MACRO PVDD2ANA
    CLASS PAD ;
    FOREIGN PVDD2ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AVDD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  20.510 184.060 26.440 190.000 ;
        RECT  12.210 0.750 17.790 2.250 ;
        RECT  5.000 78.685 25.000 86.680 ;
        RECT  12.000 184.060 18.000 190.000 ;
        RECT  3.560 184.060 9.490 190.000 ;
        LAYER M1 ;
        RECT  20.510 184.060 26.440 190.000 ;
        RECT  12.210 0.750 17.790 2.250 ;
        RECT  12.000 184.060 18.000 190.000 ;
        RECT  3.560 184.060 9.490 190.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  27.940 0.000 30.000 190.000 ;
        RECT  2.060 0.000 27.940 182.560 ;
        RECT  0.000 0.000 2.060 190.000 ;
        LAYER VIA1 ;
        RECT  20.510 184.060 26.440 190.000 ;
        RECT  12.000 184.060 18.000 190.000 ;
        RECT  3.560 184.060 9.490 190.000 ;
        LAYER M2 ;
        RECT  27.940 0.000 30.000 190.000 ;
        RECT  2.060 0.000 27.940 182.560 ;
        RECT  0.000 0.000 2.060 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVDD2ANA

MACRO PVDD2DGZ
    CLASS PAD ;
    FOREIGN PVDD2DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VDDPST
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  15.605 0.750 17.075 1.005 ;
        LAYER M1 ;
        RECT  15.605 0.750 17.075 1.005 ;
        END
    END VDDPST
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVDD2DGZ

MACRO PVDD2POC
    CLASS PAD ;
    FOREIGN PVDD2POC 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VDDPST
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  15.605 0.750 17.075 1.005 ;
        LAYER M1 ;
        RECT  15.605 0.750 17.075 1.005 ;
        END
    END VDDPST
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVDD2POC

MACRO PVSS1ANA
    CLASS PAD ;
    FOREIGN PVSS1ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AVSS
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 0.750 16.465 1.365 ;
        RECT  5.000 78.685 25.000 86.685 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  14.000 0.750 16.000 1.365 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M2 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVSS1ANA

MACRO PVSS1DGZ
    CLASS PAD ;
    FOREIGN PVSS1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  22.335 186.320 25.265 190.000 ;
        RECT  17.935 186.320 20.865 190.000 ;
        RECT  13.535 0.750 16.465 1.365 ;
        RECT  5.000 78.685 25.000 86.685 ;
        RECT  13.535 186.320 16.465 190.000 ;
        RECT  9.135 186.320 12.065 190.000 ;
        RECT  4.735 186.320 7.665 190.000 ;
        LAYER M1 ;
        RECT  22.335 186.320 25.265 190.000 ;
        RECT  17.935 186.320 20.865 190.000 ;
        RECT  14.000 0.750 16.000 1.365 ;
        RECT  13.535 186.320 16.465 190.000 ;
        RECT  9.135 186.320 12.065 190.000 ;
        RECT  4.735 186.320 7.665 190.000 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 185.820 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 185.820 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 185.820 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 185.820 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 185.820 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA1 ;
        RECT  22.335 186.320 25.265 190.000 ;
        RECT  17.935 186.320 20.865 190.000 ;
        RECT  13.535 186.320 16.465 190.000 ;
        RECT  9.135 186.320 12.065 190.000 ;
        RECT  4.735 186.320 7.665 190.000 ;
        LAYER M2 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 185.820 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 185.820 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 185.820 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 185.820 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 185.820 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA2 ;
        RECT  22.335 186.320 25.265 190.000 ;
        RECT  17.935 186.320 20.865 190.000 ;
        RECT  13.535 186.320 16.465 190.000 ;
        RECT  9.135 186.320 12.065 190.000 ;
        RECT  4.735 186.320 7.665 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVSS1DGZ

MACRO PVSS2ANA
    CLASS PAD ;
    FOREIGN PVSS2ANA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AVSS
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 0.750 16.465 1.365 ;
        RECT  5.000 78.685 25.000 86.685 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  14.000 0.750 16.000 1.365 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M2 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  3.500 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVSS2ANA

MACRO PVSS2DGZ
    CLASS PAD ;
    FOREIGN PVSS2DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  5.000 78.685 25.000 86.685 ;
        END
    END VSSPST
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M5 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M6 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  16.540 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  13.460 0.910 16.540 77.185 ;
        RECT  3.500 0.000 13.460 77.185 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVSS2DGZ

MACRO PVSS3DGZ
    CLASS PAD ;
    FOREIGN PVSS3DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 190.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M7 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M6 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M5 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M4 ;
        RECT  13.620 0.000 16.380 0.750 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M3 ;
        RECT  5.000 78.685 25.000 86.685 ;
        LAYER M2 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  5.000 78.685 25.000 86.685 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA1 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M2 ;
        RECT  25.765 0.000 30.000 190.000 ;
        RECT  21.835 0.000 25.765 183.560 ;
        RECT  21.365 0.000 21.835 190.000 ;
        RECT  17.435 0.000 21.365 183.560 ;
        RECT  16.965 0.000 17.435 190.000 ;
        RECT  13.035 0.000 16.965 183.560 ;
        RECT  12.565 0.000 13.035 190.000 ;
        RECT  8.635 0.000 12.565 183.560 ;
        RECT  8.165 0.000 8.635 190.000 ;
        RECT  4.235 0.000 8.165 183.560 ;
        RECT  0.000 0.000 4.235 190.000 ;
        LAYER VIA2 ;
        RECT  22.335 184.060 25.265 190.000 ;
        RECT  17.935 184.060 20.865 190.000 ;
        RECT  13.535 184.060 16.465 190.000 ;
        RECT  9.135 184.060 12.065 190.000 ;
        RECT  4.735 184.060 7.665 190.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 190.000 ;
        LAYER M4 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M5 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M6 ;
        RECT  16.540 0.000 30.000 190.000 ;
        RECT  13.460 0.910 16.540 190.000 ;
        RECT  0.000 0.000 13.460 190.000 ;
        LAYER M7 ;
        RECT  26.500 0.000 30.000 190.000 ;
        RECT  16.540 0.000 26.500 77.185 ;
        RECT  3.500 88.185 26.500 190.000 ;
        RECT  13.460 0.910 16.540 77.185 ;
        RECT  3.500 0.000 13.460 77.185 ;
        RECT  0.000 0.000 3.500 190.000 ;
    END
END PVSS3DGZ

END LIBRARY
